/*

 n_tap_fir.v
 --------------
 By: Augustas Jackevic
 Date: February 2021

 Module Description:
 -------------------
 This module is a design of an n-type FIR (Finite Impulse Response)
 filter. This filter is the convolution operation between the
 input data (data_in) and the coefficient data (coefficient_in). The
 default LENGTH is 10. It should be noted, to help understand the workings
 of the FIR_MAIN state, the PDF in:
 The workings of an FIR filter\The workings of a FIR filter.pdf should be read.

*/

module n_tap_fir #(
	parameter LENGTH = 10,
	parameter DATA_WIDTH = 8
)(
	input clock,
	input load_coefficients_flag,
	input load_data_flag,
	input stop_data_load_flag,
	input signed [DATA_WIDTH - 1:0] coefficient_in,
	input signed [DATA_WIDTH - 1:0] data_in,
	output reg signed [18:0] data_out
);



// Creating the internal buffers for the coefficients and data in,
reg signed [DATA_WIDTH - 1:0] coeff_buffer [0:LENGTH - 1];
reg signed [DATA_WIDTH - 1:0] input_data_buffer [0:LENGTH -1];

// Coefficient counter. Filter will only for 1023 ((2^10)-1) taps.
reg [9:0] coeff_counter;

// Local parameter to store the FIR filters output.
// FIR output width = input data width + coefficient width + log2(LENGTH)
reg signed [18:0] fir_output;



// FSM states
reg [2:0] state;
reg [2:0] IDLE = 3'd0;
reg [2:0] LOAD_COEFFICIENTS = 3'd1;
reg [2:0] FIR_MAIN = 3'd2;
reg [2:0] STOP = 3'd3;




// Setting the initial values.
initial begin : init_values

	// Set all the values inside the coeff_buffer to 0.
	integer k;
	for (k = 0; k <= LENGTH - 1 ; k = k + 1) begin
		coeff_buffer[k] = 0;
		input_data_buffer[k] = 0;
	end

	// Set the internal variables and outputs to 0.
	state = IDLE;
	coeff_counter = 0;
	data_out = 0;
	fir_output = 0;
end





integer n;
always @(posedge clock) begin
	case(state)
	
	
		// State IDLE. This checks the load_coefficients_flag value and only
		// transition to state LOAD_COEFFICIENTS when the flag is high.
		IDLE: begin
			if(load_coefficients_flag == 1) begin
				state = LOAD_COEFFICIENTS;
			end
		end
		
		
		
		// State LOAD_COEFFICIENTS. This state is responsiable for loading the
		// coefficients to coeff_buffer. Once all the coefficients are loaded the
		// state transitions to FIR_MAIN.
		LOAD_COEFFICIENTS: begin
		
			// A for loop that shifts the values inside coeff_buffer by 1 position.
			for (n = LENGTH - 1; n > 0; n = n - 1) begin
				coeff_buffer[n] <= coeff_buffer[n-1];
			end

			// Load the new coefficient value to the start of coeff_buffer.
			coeff_buffer[0] <= coefficient_in;

			// Increment coeff_counter, when it is equal to LENGTH, the
			// coeff_buffer is full, thus transition to state FIR_MAIN.
			coeff_counter = coeff_counter + 10'd1;
			if(coeff_counter == LENGTH) begin
				state = FIR_MAIN;
			end
		end
		
		
		// State FIR_MAIN. This state is responsiable for the main FIR opperation. It follows
		// the logic outlined in the pdf "The workings of a FIR filter".
		FIR_MAIN: begin
		
			// If the data input stream is ready, do the following.
			if(load_data_flag == 1) begin
				//Shift the values inside input_data_buffer by 1.
				for (n = LENGTH - 1; n > 0; n = n - 1) begin
					input_data_buffer[n] <= input_data_buffer[n - 1];
				end

				// Load the new data_in value to the start of input_data_buffer.
				input_data_buffer[0] <= data_in;
			
				// fir_output is set to 0, as everytime FIR_MAIN loops, previous fir_output value is used, hence the first
				// fir_output value that is used in the for loop would not be of the correct value.
				fir_output = 0;
				// A multiplication between the input data and the corresponding coefficients
				// in the delayed buffer line. This for loop also sums all the components together.
				for (n = 0; n <= LENGTH - 1; n = n + 1) begin
					fir_output = fir_output + (input_data_buffer[n] * coeff_buffer[LENGTH - 1 - n]);
				end
			end

			// Load the output of the FIR to the output reg of the module, data_out.
			data_out = fir_output;
			
			// Transition to stop state when stop_data_load_flag is 1.
			if(stop_data_load_flag == 1) begin
				state = STOP;
			end
		end

		
		STOP: begin

		end
		
		// State default. This state is added just incase the FSM is in an unknown state, it resets all
		// all the local parameter and sets state to IDLE.
		default: begin
			// Set all the values inside the coeff_buffer to 0.
			integer k;
			for (k = 0; k <= LENGTH - 1 ; k = k + 1) begin
				coeff_buffer[k] = 0;
				input_data_buffer[k] = 0;
			end

			// Set the internal variables and outputs to 0.
			state = IDLE;
			coeff_counter = 0;
			data_out = 0;
			fir_output = 0;
		end

	endcase

end



endmodule
