module testMIFRead #(
	parameter LENGTH = 20000,
	parameter DATA_WIDTH = 13

)(
	input clock,
	input enable,
	
	output reg signed [DATA_WIDTH - 1:0] outputValue
);




endmodule
