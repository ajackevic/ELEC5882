module squareRootCal(
	
);


endmodule
