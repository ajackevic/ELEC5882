module testMIFRead(


);




endmodule
