module absolute_value_tb;



endmodule
