/*

 matched_filter.v
 --------------
 By: Augustas Jackevic
 Date: July 2021

 Module Description:
 -------------------
 This module creates the matched filter. The matched filter is the convelution opperation
 between the input data and the matched filter impulse response (very over-simplifyied). Both
 signals are applied through a hilbert transform filter (removed the negative frequencies) and then
 conveluted. The hilbert transform is required to avoide alliasying. Due to the hiolbert transform, a
 complex signal is aquired thus a comple FIR filter is utalised for the convelution.
 
 In this module, the matched filter coefficients are aquired from the MFImpulseCoeff MIF file (coefficients
 are obtained from MATLAB), and the input data is read from the MFInputData MIF file. This data is then applied
 through the hilbert transform module to aquire a complex signal. The coefficients are loaded to the complex
 FIR filter and the data in complex signal is then applied to the FIR filter, with the output being the convelution
 product between the matched filter impulse response coefficients and the applied data in.


*/


module matched_filter #(
	parameter COEFF_LENGTH = 10000,
	parameter DATA_LENGTH = 330000,
	parameter HT_COEFF_LENGTH = 27,
	parameter HT_DATA_WIDTH = 18,
	parameter DATA_WIDTH = 18
)(
	input clock,
	input enable,
	
	output reg signed [DATA_WIDTH - 1:0] filterOut  // This will need to be *3 ot *4?
);


// Local parameters for the module read_MIF_file.
localparam COEFF = 1;
localparam DATA_IN = 2;


// Enable regs for the instantiated modules.
reg enableMFCoeff;
reg enableMFDataIn;
reg enablecomplexFIRCoeff;
reg enableHT;
reg enableComplexFIRData;


// A reg for informing the complex FIR filter when the data is about to be stopped.
reg stopDataLoadFlag;


// Output ports for the instantiated modules.
wire coeffFinishedFlag;
wire dataInFinishedFlag;
wire signed [DATA_WIDTH - 1:0] coeffMIFOutRe;
wire signed [DATA_WIDTH - 1:0] coeffMIFOutIm;
wire signed [DATA_WIDTH - 1:0] dataMIFOutRe;

wire signed [(DATA_WIDTH * 2) - 1:0] HTOutRe;
wire signed [(DATA_WIDTH * 2) - 1:0] HTOutIm;

wire signed [(DATA_WIDTH * 3) - 1:0] MFOutputRe;
wire signed [(DATA_WIDTH * 3) - 1:0] MFOutputIm;



// FSM
reg [2:0] state;
localparam IDLE = 1;
localparam LOAD_COEFF = 2;
localparam LOAD_DATA = 3;
localparam STOP = 4;




// Set the initial values of the local parameters.
initial begin

	enableMFCoeff <= 1'd0;
	enableMFDataIn <= 1'd0;
	enablecomplexFIRCoeff <= 1'd0;
	enableHT <= 1'd0;
	
	
	enableComplexFIRData <= 1'd0;
	stopDataLoadFlag <= 1'd0;
	
	
	state <= IDLE;
	filterOut <= {(DATA_WIDTH){1'd0}};
end




// Instantiating the module read_MIF_file. This is used to read the coefficients from the MFImpulseCoeff.mif file.
read_MIF_file #(
	.LENGTH 				(COEFF_LENGTH),
	.DATA_WIDTH 		(DATA_WIDTH),
	.DATA_TYPE 			(COEFF)

) MFCoeff (
	.clock				(clock),
	.enable				(enableMFCoeff),
	
	.dataFinishedFlag	(coeffFinishedFlag),	
	.outputRe			(coeffMIFOutRe),
	.outputIm			(coeffMIFOutIm)
);




// Instantiating the module read_MIF_file. This is used to read the data in from the MFInputData.mif file. 
read_MIF_file #(
	.LENGTH 				(DATA_LENGTH),
	.DATA_WIDTH 		(DATA_WIDTH),
	.DATA_TYPE 			(DATA_IN)

) MFDataIn (
	.clock				(clock),
	.enable				(enableMFDataIn),
	
	.dataFinishedFlag	(dataInFinishedFlag),	
	.outputRe			(dataMIFOutRe),
	.outputIm			()
);





// Instantiating the module n_tap_complex_fir. This is used for the main opperation of the matched filter
// between the complex input data and the complex impulse reponse of the matched filter.
n_tap_complex_fir #(
	.LENGTH					(COEFF_LENGTH * 2),
	.DATA_WIDTH 			(DATA_WIDTH)
) coplexFIR (
	.clock					(clock),
	.loadCoeff				(enablecomplexFIRCoeff),
	.coeffSetFlag			(coeffFinishedFlag),
	.loadDataFlag			(enableComplexFIRData),
	.stopDataLoadFlag		(stopDataLoadFlag),
	.dataInRe				(HTOutRe),
	.dataInIm				(HTOutIm),
	.coeffInRe				(coeffMIFOutRe),
	.coeffInIm				(coeffMIFOutIm),
	
	.dataOutRe				(MFOutputRe),
	.dataOutIm				(MFOutputIm)
);





// Instantiating the module hilbert_transform. This is used to aquire a complex signal from a real signal 
// by performing hilbert transform filtering of the data aquired from MFInputData.mif.
 hilbert_transform #(
	.LENGTH 				(HT_COEFF_LENGTH),
	.DATA_WIDTH 		(DATA_WIDTH)
) hilbertTransform (
	.clock				(clock),
	.enable				(enableHT),
	.stopDataInFlag	(),
	.dataIn				(dataMIFOutRe),
	
	.dataOutRe			(HTOutRe),
	.dataOutIm			(HTOutIm)
);







always @ (posedge clock) begin
	case(state)
		
		// State IDLE. This state waits until enable is set before transistioning to LOAD_COEFF.
		IDLE: begin
			if(enable) begin
				state <= LOAD_COEFF;
			end
			else begin
				filterOut <= {(DATA_WIDTH){1'd0}}; // This will need to be *3 ot *4?
			end
		end
		
		
		// State LOAD_COEFF. This state enables the majority of the enable regs for the instantiated modules.
		LOAD_COEFF: begin
						
			if(coeffFinishedFlag) begin
			
				enableMFCoeff <= 1'd0;
				state <= LOAD_DATA;
				enableMFDataIn <= 1'd1;
				enableHT <= 1'd1;
				
			end
			else begin
				enableMFCoeff <= 1'd1;
				enableMFDataIn <= 1'd1;
				enablecomplexFIRCoeff <= 1'd1;
				enableHT <= 1'd1;
				enableComplexFIRData <= 1'd1;
			end
		end
		
		LOAD_DATA: begin
		
		end
		
		STOP: begin
		
		end
		
		default: begin
		
		end
		
	endcase
end

/*
 Right in this script I need to instantiate the n_tap_complex_fir module and setup_MF_coeff.
 I then need to pass on coefficient values from setup_MF_coeff to n_tap_complex_fir. Then I 
 need edit the script setup_MF_coeff so that its compatiable with two types of MIF file
 (have it based on pre set parameters). Hence that module can be used to read two MIF files,
 thus will need two instantiations. Once the coefficients are set (could potentially be done 
 in parallel), send through the x_t data to n_tap_complex_fir. The output should then go 
 through an ABS algorithm (obtains the absloute value of y_t).
*/

endmodule
