module  absolute_value(


);


endmodule
