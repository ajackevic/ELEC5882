module testMIFRead_tb;




endmodule
