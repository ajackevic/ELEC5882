module matched_filter_tb;


endmodule
