module matched_filter(


);



endmodule
