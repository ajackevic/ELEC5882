module squareRootCal_tb;



endmodule;
