module hilbert_transform_tb;


endmodule
