module setupComplexCoefficients)(


);



endmodule
