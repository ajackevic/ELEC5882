module setup_HT_coeff


endmodule
