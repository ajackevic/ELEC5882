module setup_complex_coefficients_tb;



endmodule
